library ieee;
use ieee.std_logic_1164.all;

entity bus_interface_cu is
  port (RESET, CLOCK                                               : in  std_logic;
        CS_cu, R_Wn_cu                                             : in  std_logic;
        EN_STATE                                                   : out std_logic_vector (2 downto 0);
        ADD_cu                                                     : in  std_logic_vector (2 downto 0);
        SEL_mux_cu, ATN_cu, EN_regCTRL, EN_regDATARX, EN_regDATATX : out std_logic;
        TX_ack_cu                                                  : out std_logic;
        RX_ack_cu                                                  : out std_logic;
        CLRatn_cu                                                  : in  std_logic;
        RX_FULL_cu, TX_EMPTY_cu, ERROR_cu, ATNack_cu               : in  std_logic);
end bus_interface_cu;


architecture behav of bus_interface_cu is


  type state_type is (IDLE,
                      WRITE_CTRL,
                      WAIT_s,
                      WRITE_CTRL_ATN,
                      READ_STATUS,
                      WRITE_TXdata,
                      READ_RXdata,
                      ATN_TX_s,
                      ATN_RX_or_ERROR_s,
                      ATN_TXand_RX_or_ERROR_s,
                      ATN_OVERRUN_s,
                      ATN_OVERRUNandTX_s,
                      CLEAR_s
                      );

  signal present_state : state_type;

begin
  state_update : process(CLOCK, RESET)
  begin
    if (RESET = '0') then
      present_state <= IDLE;

    elsif (CLOCK'event and CLOCK = '1') then

      case present_state is

        when IDLE =>
          if((TX_EMPTY_cu = '1') and (RX_FULL_cu = '1') and (ERROR_cu = '1')) then present_state  <= ATN_OVERRUNandTX_S;
          elsif (TX_EMPTY_cu = '1') and ((RX_FULL_cu = '1' or ERROR_cu = '1')) then present_state <= ATN_TXand_RX_or_ERROR_s;
          elsif (RX_FULL_cu = '1') and(ERROR_cu = '1') then present_state                         <= ATN_OVERRUN_s;
          elsif (TX_EMPTY_cu = '1') then present_state                                            <= ATN_TX_s;
          elsif (RX_FULL_cu = '1' or ERROR_cu = '1') then present_state                           <= ATN_RX_or_ERROR_s;

          elsif (CS_cu = '1' and R_Wn_cu = '0' and ADD_cu = "011") then present_state <= WRITE_CTRL;
          else present_state                                                          <= IDLE;
          end if;

        when WRITE_CTRL =>
          if (CS_cu = '1' and R_Wn_cu = '1' and ADD_cu = "010") then present_state    <= READ_STATUS;
          elsif (CS_cu = '1' and R_Wn_cu = '0' and ADD_cu = "000") then present_state <= WRITE_TXdata;
          else present_state                                                          <= WAIT_s;
--per gestire ritardo nella risposta tra tx e bus
          end if;

        when WAIT_s => present_state <= IDLE;


        when READ_STATUS =>
          if (RX_FULL_cu = '1' and CS_cu = '1' and R_Wn_cu = '1' and ADD_cu = "001") then present_state     <= READ_RXdata;
          elsif (TX_EMPTY_cu = '1' and CS_cu = '1' and R_Wn_cu = '0' and ADD_cu = "000") then present_state <= WRITE_TXdata;
          elsif (CS_cu = '1' and R_Wn_cu = '0' and ADD_cu = "011") then present_state                       <= WRITE_CTRL;
          elsif (CS_cu = '1' and R_Wn_cu = '1' and ADD_cu = "010") then present_state                       <= READ_STATUS;
          else present_state                                                                                <= IDLE;
          end if;


        when WRITE_TXdata =>
          present_state <= IDLE;

        when READ_RXdata =>
          if(TX_EMPTY_cu = '1' and CS_cu = '1' and R_Wn_cu = '0' and ADD_cu = "000") then present_state <= WRITE_TXdata;
          else present_state                                                                            <= IDLE;
          end if;

        when WRITE_CTRL_ATN => present_state <= CLEAR_s;

        when CLEAR_s =>
          if (CS_cu = '1' and R_Wn_cu = '1' and ADD_cu = "010") then present_state <= READ_STATUS;
          else present_state                                                       <= IDLE;
          end if;

        when ATN_TX_s =>
          if (RX_FULL_cu = '1') and (ERROR_cu = '1') then present_state               <= ATN_OVERRUNandTX_s;
          elsif (RX_FULL_cu = '1' or ERROR_cu = '1') then present_state               <= ATN_TXand_RX_or_ERROR_s;
          elsif (CLRatn_cu = '1' or ATNack_cu = '1') then present_state               <= CLEAR_s;
          elsif (CS_cu = '1' and R_Wn_cu = '0' and ADD_cu = "011") then present_state <= WRITE_CTRL_ATN;
          else present_state                                                          <= ATN_TX_s;
          end if;

        when ATN_RX_or_ERROR_S =>
          if (TX_EMPTY_cu = '1' and ERROR_cu = '1' and RX_FULL_cu = '1') then present_state <= ATN_OVERRUNandTX_s;
          elsif (TX_EMPTY_cu = '1') then present_state                                      <= ATN_TXand_RX_or_ERROR_s;
          elsif (RX_FULL_cu = '1' and ERROR_cu = '1') then present_state                    <= ATN_OVERRUN_s;
          elsif (CLRatn_cu = '1' or ATNack_cu = '1') then present_state                     <= CLEAR_s;
          elsif (CS_cu = '1' and R_Wn_cu = '0' and ADD_cu = "011") then present_state       <= WRITE_CTRL_ATN;
          else present_state                                                                <= ATN_RX_or_ERROR_s;
          end if;

        when ATN_TXand_RX_or_ERROR_s =>
          if (TX_EMPTY_cu = '1' and RX_FULL_cu = '1' and ERROR_cu = '1') then present_state <= ATN_OVERRUNandTX_s;
          elsif (CLRatn_cu = '1' or ATNack_cu = '1') then present_state                     <= CLEAR_s;
          elsif (CS_cu = '1' and R_Wn_cu = '0' and ADD_cu = "011") then present_state       <= WRITE_CTRL_ATN;
          else present_state                                                                <= ATN_TXand_RX_or_ERROR_s;
          end if;

        when ATN_OVERRUN_s =>
          if (TX_EMPTY_cu = '1') then present_state                                   <= ATN_OVERRUNandTX_s;
          elsif (CLRatn_cu = '1' or ATNack_cu = '1') then present_state               <= CLEAR_s;
          elsif (CS_cu = '1' and R_Wn_cu = '0' and ADD_cu = "011") then present_state <= WRITE_CTRL_ATN;
          else present_state                                                          <= ATN_OVERRUN_s;
          end if;

        when ATN_OVERRUNandTX_s =>
          if (CLRatn_cu = '1' or ATNack_cu = '1') then present_state                  <= CLEAR_s;
          elsif (CS_cu = '1' and R_Wn_cu = '0' and ADD_cu = "011") then present_state <= WRITE_CTRL_ATN;
          else present_state                                                          <= ATN_OVERRUNandTX_s;
          end if;

        when others =>
          present_state <= IDLE;
      end case;
    end if;
  end process;


  FSM_cu : process(present_state)
  begin



    --default values

    SEL_mux_cu   <= '1';  --LO LASCIO DI DEFAULT A ZERO COSI DA POTER MANDARE SEMPRE L'ERRORE SU DOUT
    EN_regCTRL   <= '0';
    EN_regDATARX <= '0';
    EN_regDATATX <= '0';
    TX_ack_cu    <= '0';
    EN_regDATARX <= '0';
    EN_STATE(0)  <= '1';
    EN_STATE(1)  <= '1';
    EN_STATE(2)  <= '1';  --LO LASCIO SEMPRE ALTO COSI DA POTER SEMPRE SENTIRE L'ERRORE
    ATN_cu       <= '0';
    RX_ack_cu    <= '0';

    case present_state is
      when IDLE =>
        SEL_mux_cu <= '1';
        ATN_cu     <= '0';

      when WRITE_CTRL =>
        EN_regCTRL <= '1';
        ATN_cu     <= '0';

      when WAIT_s =>
        ATN_cu <= '0';

      when WRITE_CTRL_ATN =>
        EN_regCTRL  <= '1';
        ATN_cu      <= '1';
        EN_STATE(0) <= '0';
        EN_STATE(1) <= '0';
        EN_STATE(2) <= '0';

      when READ_STATUS =>
        SEL_MUX_cu  <= '1';
        ATN_cu      <= '0';
        EN_STATE(0) <= '0';
        EN_STATE(1) <= '0';
        EN_STATE(2) <= '0';

      when READ_RXdata =>               -- LEGGO RX_DATA
        SEL_mux_cu   <= '0';
        EN_regDATARX <= '1';
        ATN_cu       <= '0';
        RX_ack_cu    <= '1';
        TX_ack_cu    <= '0';

      when WRITE_TXdata =>              -- SCRIVO SU TX_DATA
        EN_regDATATX <= '1';
        ATN_cu       <= '0';
        TX_ack_cu    <= '1';

      when ATN_TX_s =>
        ATN_cu      <= '1';
        EN_STATE(0) <= '1';
        EN_STATE(1) <= '0';
        EN_STATE(2) <= '1';
        SEL_MUX_cu  <= '1';

      when ATN_RX_or_ERROR_s =>
        ATN_cu       <= '1';
        EN_regDATARX <= '1';
        EN_STATE(0)  <= '0';
        EN_STATE(1)  <= '1';
        EN_STATE(2)  <= '0';
        SEL_MUX_cu   <= '1';

      when ATN_TXand_RX_or_ERROR_s =>
        ATN_cu       <= '1';
        EN_regDATARX <= '1';
        EN_STATE(0)  <= '0';
        EN_STATE(1)  <= '0';
        EN_STATE(2)  <= '0';
        SEL_MUX_cu   <= '1';

      when ATN_OVERRUN_s =>
        ATN_cu      <= '1';
        EN_STATE(0) <= '0';
        EN_STATE(1) <= '1';
        EN_STATE(2) <= '0';
        SEL_MUX_cu  <= '1';

      when ATN_OVERRUNandTX_s =>
        ATN_cu      <= '1';
        EN_STATE(0) <= '0';
        EN_STATE(1) <= '0';
        EN_STATE(2) <= '0';
        SEL_MUX_cu  <= '1';


      when CLEAR_s =>
        ATN_cu      <= '0';
        EN_STATE(0) <= '0';
        EN_STATE(1) <= '0';
        EN_STATE(2) <= '0';




    end case;
  end process;

end behav;
