-------------------------------------------------------------------------------
-- Title      : UART
-- Project    : 
-------------------------------------------------------------------------------
-- File       : uart.vhd
-- Author     : wackoz  <wackoz@wT14s>
-- Company    : 
-- Created    : 2021-01-07
-- Last update: 2021-02-02
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: UART
-------------------------------------------------------------------------------
-- Copyright (c) 2021 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2021-01-07  1.0      wackoz  Created
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- Title      : Uart
-- Project    : UART
-------------------------------------------------------------------------------
-- File       : uart.vhd


library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity uart is

  port (
    clock  : in  std_logic;
    reset  : in  std_logic;
    RxD    : in  std_logic;
    TxD    : out std_logic;
    Dout   : out std_logic_vector(7 downto 0);
    Din    : in  std_logic_vector(7 downto 0);
    ATN    : out std_logic;
    ATNACK : in  std_logic;
    ADD    : in  std_logic_vector(2 downto 0);
    R_Wn   : in  std_logic;
    CS     : in  std_logic
    );

end uart;

-------------------------------------------------------------------------------

architecture str of uart is

  -----------------------------------------------------------------------------
  -- Internal signal declarations
  -----------------------------------------------------------------------------

  signal p_in          : std_logic_vector(7 downto 0);
  signal tx_empty_ack  : std_logic;
  signal status_rx_full       : std_logic;
  signal status_flag_error    : std_logic;
  signal Pout          : std_logic_vector(7 downto 0);
  signal TX_out        : std_logic_vector(7 downto 0);
  signal RX_in         : std_logic_vector(7 downto 0);
  signal tx_empty      : std_logic;
  signal TX_ACK        : std_logic;
  signal RX_ACK        : std_logic;
  signal RX_ENABLE     : std_logic;
  signal TX_ENABLE     : std_logic;
  signal CLRatn        : std_logic;
  signal SEL_MUX       : std_logic;
  signal FF_IN         : std_logic_vector(2 downto 0);
  signal FF_OUT        : std_logic_vector(2 downto 0);
  signal ENABLE_FF     : std_logic_vector(2 downto 0);
  signal FF_IN_tmp     : std_logic_vector(2 downto 0);
  signal rx_enable_tmp : std_logic;


  component tx is
    port (
      clock        : in  std_logic;
      reset        : in  std_logic;
      tx_enable    : in  std_logic;
      p_in         : in  std_logic_vector(7 downto 0);
      TxD          : out std_logic;
      tx_empty     : out std_logic;
      tx_empty_ack : in  std_logic);
  end component tx;



  component rx is
    port (
      clock      : in  std_logic;
      reset      : in  std_logic;
      rx_enable  : in  std_logic;
      rx_ack     : in  std_logic;
      rxD        : in  std_logic;
      status_rx_full    : out std_logic;
      status_flag_error : out std_logic;
      Pout       : out std_logic_vector(7 downto 0));
  end component rx;

  component BUS_INTERFACE is
    port (
      Dout                 : out std_logic_vector (7 downto 0);
      TX_out               : out std_logic_vector (7 downto 0);
      RX_in, Din           : in  std_logic_vector (7 downto 0);
      CLOCK, RESET         : in  std_logic;
      RX_ENABLE, TX_ENABLE : out std_logic;
      ATNack               : in  std_logic;
      ATN, TX_ACK, RX_ACK  : out std_logic;
      FF_IN_B              : in  std_logic_vector (2 downto 0);
      ADD                  : in  std_logic_vector (2 downto 0);
      R_Wn, CS             : in  std_logic);
  end component BUS_INTERFACE;


begin

  trasmettitore : tx port map (
    clock        => clock,
    reset        => reset,
    tx_enable    => TX_ENABLE,
    p_in         => TX_out,
    tx_empty_ack => TX_ACK,             --vedi bene
    tx_empty     => tx_empty,
    TxD          => TxD);

  ricevitore : rx port map (
    clock      => clock,
    reset      => reset,
    rx_enable  => RX_ENABLE,
    rx_ack     => rx_ack,
    rxD        => RxD,
    status_rx_full    => status_rx_full,
    status_flag_error => status_flag_error,
    Pout       => Pout);


  -- instance "BUS_INTERFACE_1"
  BUS_INTERFACE_1 : BUS_INTERFACE
    port map (
      Dout      => Dout,
      TX_out    => TX_out,
      RX_in     => Pout,
      Din       => Din,
      CLOCK     => CLOCK,
      RESET     => RESET,
      RX_ENABLE => RX_ENABLE,
      TX_ENABLE => TX_ENABLE,
      ATNack    => ATNack,
      ATN       => ATN,
      TX_ACK    => TX_ACK,
      rx_ack    => rx_ack,
      FF_IN_B   => FF_IN_tmp,
      ADD       => ADD,
      R_Wn      => R_Wn,
      CS        => CS);

  FF_IN_tmp <= (status_flag_error)&(tx_empty)&(status_rx_full);



end architecture str;

-------------------------------------------------------------------------------
