-------------------------------------------------------------------------------
-- Title      : Testbench for design "uart"
-- Project    : 
-------------------------------------------------------------------------------
-- File       : uart_tb.vhd
-- Author     : wackoz  <wackoz@wT14s>
-- Company    : 
-- Created    : 2021-01-07
-- Last update: 2021-02-06
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2021 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2021-01-07  1.0      wackoz  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity uart_tb is

end entity uart_tb;

-------------------------------------------------------------------------------

architecture arch of uart_tb is

  -- component ports
  signal clock  : std_logic := '1';
  signal reset  : std_logic;
  signal RxD    : std_logic;
  signal TxD    : std_logic;
  signal Dout   : std_logic_vector(7 downto 0);
  signal Din    : std_logic_vector(7 downto 0);
  signal ATN    : std_logic;
  signal ATNACK : std_logic;
  signal ADD    : std_logic_vector(2 downto 0);
  signal R_Wn   : std_logic;
  signal CS     : std_logic;


begin  -- architecture arch

  -- component instantiation
  DUT : entity work.uart
    port map (
      clock  => clock,
      reset  => reset,
      RxD    => RxD,
      TxD    => TxD,
      Dout   => Dout,
      Din    => Din,
      ATN    => ATN,
      ATNACK => ATNACK,
      ADD    => ADD,
      R_Wn   => R_Wn,
      CS     => CS);

  -- clock generation
  clock <= not clock after 31.25 ns;

  -- waveform generation
  WaveGen_Proc : process
  begin
    reset <= '0';
    ADD <="000";
    R_Wn <= '0';
    CS <= '0';
    Din <= "00000000";
    ATNack<='0';
    wait for 62.5 ns;
    reset <= '1';
    ADD   <= "011";  -- VADO A SCRIVERE NEL REG DI CONTROLLO
    R_Wn  <= '0';
    CS    <= '1';
    wait for 62.5 ns;
    Din <= "00000010";
    ADD   <= "000";
    R_Wn  <= '0';
    wait for 62.5 ns;
    Din   <= "10011000";   -- trasmetto la parola a TXDATA
    wait for 62.5 ns;
    ADD   <= "010";   --leggo lo stato
    R_Wn  <= '1';
    wait for 62.5 ns;
    CS <= '0';
    ADD <="000";
    wait for 86.875 us;
    ATNack <= '1';
    wait for 62.5 ns;
    ADD  <= "010";
    CS   <= '1';
    R_Wn <= '1';  --leggo lo stato e controllo se rxfull � alto e se il
    --trasmettitore ha concluso la trasmissione
    wait for 62.5 ns;
    ATNACK <='0';
    ADD <= "011";    --ABILITO RX e spengo TX
    CS <= '1';
    R_Wn <= '0';
    wait for 62.5 ns;
    Din <= "00000001";
    CS <= '0';
    ADD <="000";
    wait for 62.5 ns;
    --affronto il caso in cui sia avvenuta una ricezione corretta
    rxd <= '0';                         --
    wait for 8.6956 us;
    rxd <= '1';                         -- D0
    wait for 8.6956 us;
    rxd <= '0';                         -- D1
    wait for 8.6956 us;
    rxd <= '0';                         --D2
    wait for 8.6956 us;
    rxd <= '1';                         --D3
    wait for 8.6956 us;
    rxd <= '0';                         --D4
    wait for 8.6956 us;
    rxd <= '1';                         --D5
    wait for 8.6956 us;
    rxd <= '0';                         --D6
    wait for 8.6956 us;
    rxd <= '0';                         --D7
    wait for 8.6956 us;
    rxd <= '1';                         --corretta
    wait for 8.9456 us; --tempo necessario per trasmettere ultimo simbolo(139Tclk)+t
                        --di delay(3Tclk)+tempo di risposta esterno(1Tclk)
    CS <='1';
    ATNack <= '1';
    wait for 62.5 ns;
    ATNack <= '0';
    ADD  <= "010";
    R_Wn <= '1';  --leggo lo stato e controllo se rxfull � alto
    wait for 62.5 ns;
    ADD <= "001";
    wait for 62.5 ns; -- parola ricevuta in uscita READ_RXDATA
    --spengo ricevitore e trasmettitore
    ADD  <= "011";
    CS   <= '1';
    R_Wn <= '0';
    Din  <= "00000001";
    wait for 62.5 ns;
    ADD  <= "011";
    CS   <= '1';
    R_Wn <= '0';
    Din  <= "00000000";
    wait for 62.5 ns;
    CS <= '0';
    wait;



  end process WaveGen_Proc;

end architecture arch;

-------------------------------------------------------------------------------

configuration uart_tb_arch_cfg of uart_tb is
  for arch
  end for;
end uart_tb_arch_cfg;

-------------------------------------------------------------------------------
