library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity butterfly is
  port (
    clock
  ) ;
end butterfly ; 

architecture myArch of butterfly is

begin

end architecture ;