library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controlunit_butterfly is

  port (start             : in  std_logic;
        clock, reset      : in  std_logic;
        datapath_commands : out std_logic_vector (15 downto 0);
        done              : out std_logic);
end controlunit_butterfly;

-------------------------------------------------------------------------------

architecture behav of controlunit_butterfly is

  -----------------------------------------------------------------------------
  -- COMPONENTS
  -----------------------------------------------------------------------------

  component microROM is

    generic (constant N : integer := 24);
    port (ADDRESS                   : in  std_logic_vector (3 downto 0);
          OUT_MEM_even, OUT_MEM_odd : out std_logic_vector (N-1 downto 0));
  end component;

  component PLA_status is
    port (start, lsb_in : in  std_logic;
          cc_validation : in  std_logic_vector(1 downto 0);
          LSB_out       : out std_logic);
  end component;

  component reg is
    generic (
      N : integer);
    port (
      D                    : in  std_logic_vector(N-1 downto 0);
      clock, reset, enable : in  std_logic;
      Q                    : out std_logic_vector(N-1 downto 0));
  end component reg;

  component reg_neg_triggered is
    generic (
      N : integer);
    port (
      D                    : in  std_logic_vector(N-1 downto 0);
      clock, reset, enable : in  std_logic;
      Q                    : out std_logic_vector(N-1 downto 0));
  end component reg_neg_triggered;

  -----------------------------------------------------------------------------
  -- SIGNALS
  -----------------------------------------------------------------------------

  signal mem_out1, mem_out2, mux_out, out_uIR : std_logic_vector (23 downto 0);
  signal in_uAR_LSB                      : std_logic;
  signal out_uAR, D_uAR                       : std_logic_vector(4 downto 0);
  signal in_uAR_ADD                              : std_logic_vector(3 downto 0);

-------------------------------------------------------------------------------
begin

  --microIR fields:
  datapath_commands <= out_uIR(20 downto 5);
  done              <= out_uIR(21);
  in_uAR_ADD        <= out_uIR(4 downto 1);
  D_uAR             <= in_uAr_ADD & in_uAR_LSB;


  --instance microROM
  microROM_inst : microROM
    port map (ADDRESS      => out_uAR(4 downto 1),
              OUT_MEM_even => mem_out1,
              OUT_MEM_odd  => mem_out2);


  mux2_to_1_microROM : process(mem_out1, mem_out2, out_uAR(0)) is
  begin  -- process mux2_to_1_microROM
    if out_uAR(0) = '1' then
      mux_out <= mem_out2;
    else
      mux_out <= mem_out1;
    end if;
  end process mux2_to_1_microROM;

  --instance "late_status"
  late_status : PLA_status
    port map (start         => start,
              lsb_in        => out_uIR(0),
              cc_validation => out_uIR(23 downto 22),
              LSB_out       => in_uAR_LSB);


  -- instance "reg_uAR"
  reg_uAR : reg_neg_triggered
    generic map (
      N => 5)
    port map (
      D      => D_uAR,
      clock  => clock,
      reset  => reset,
      enable => '1',
      Q      => out_uAR);

  -- instance "reg_uIR"
  reg_uIR : reg
    generic map (
      N => 24)
    port map (
      D      => mux_out,
      clock  => clock,
      reset  => reset,
      enable => '1',
      Q      => out_uIR);



end behav;

