library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity butterfly_tb is

end entity butterfly_tb;

-------------------------------------------------------------------------------

architecture arch of butterfly_tb is

  -- component ports
  signal start,full_speed ,done                            : std_logic;
  signal AR,AI,BR,BI,WR,WI                          : std_logic_vector (19 downto 0);
  signal AR_out,AI_out,BR_out,BI_out                              : std_logic_vector (19 downto 0);

  -- clock
  signal clock : std_logic := '1';

begin  -- architecture arch

  -- component instantiation
  DUT : entity work.butterfly
    port map (
	 clock => clock,
      start => start,
		full_speed => full_speed,
		done => done,
		AR => AR,
		AI => AI,
		BR => BR,
		BI => BI,
		WR => WR,
		WI => WI,
		AR_out => AR_out,
		AI_out => AI_out,
		BR_out => BR_out,
		BI_out => BI_out
     );

  -- clock generation
  clock <= not clock after 10 ns;

  -- waveform generation
  WaveGen_Proc : process
  begin
    -- insert signal assignments here


start <= '0';
full_speed <= '0';
wait for 50 ns;
start <= '0';
full_speed <= '0';
WR <= "00000000000000000001";
WI <= "00000000001000000000";
AR <= "00000000000000000001";
AI <= "00000000001000000000";
BR <= "00000000000000000001";
BI <= "00000000001000000000";

wait for 50 ns;
start <= '1';
full_speed <= '0';
WR <= "00000000000000000001";
WI <= "00000000001000000000";
AR <= "00000000000000000001";
AI <= "00000000001000000000";
BR <= "00000000000000000001";
BI <= "00000000001000000000";
wait for 50 ns;
start <= '1';
full_speed <= '0';
WR <= "00000000000000000001";
WI <= "00000000001000000000";
AR <= "00000000000000000001";
AI <= "00000000001000000000";
BR <= "00000000000000000001";
BI <= "00000000001000000000";
wait for 50 ns;

start <= '0';
full_speed <= '0';
WR <= "00000000000000000001";
WI <= "00000000001000000000";
AR <= "00000000000000000001";
AI <= "00000000001000000000";
BR <= "00000000000000000001";
BI <= "00000000001000000000";
wait;
  end process WaveGen_Proc;



end architecture arch;