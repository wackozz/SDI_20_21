-------------------------------------------------------------------------------
-- Title      : adder
-- Project    : 
-------------------------------------------------------------------------------
-- File       : adder.vhd
-- Author     : wackoz  <wackoz@wT14s>
-- Company    : 
-- Created    : 2020-12-26
-- Last update: 2021-01-09
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: adder/subtractor Nbit
-------------------------------------------------------------------------------
-- Copyright (c) 2020 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2020-12-26  1.0      wackoz  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-------------------------------------------------------------------------------

entity adder is

  generic (
    N : integer := 4);

  port (
    clock   : in  std_logic;
    reset   : in  std_logic;
    add_sub : in  std_logic;
    A       : in  std_logic_vector(N-1 downto 0);
    B       : in  std_logic_vector(N-1 downto 0);
    Y       : out std_logic_vector(N downto 0));

end entity adder;

-------------------------------------------------------------------------------

architecture str of adder is
begin
  sum : process (clock, reset) is
  begin  -- process sum
    if reset = '0' then                     -- asynchronous reset (active low)
      Y <= (others => '0');
    elsif clock'event and clock = '1' then  -- rising clock edge
      if(add_sub = '0') then
        Y <= std_logic_vector(resize(signed(A), N+1)+resize(signed(B), N+1));
      else
        Y <= std_logic_vector(resize(signed(A), N+1)-resize(signed(B), N+1));
      end if;
    end if;
  end process sum;
end architecture str;

-------------------------------------------------------------------------------
